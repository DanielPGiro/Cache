--
-- Entity: negative edge triggered 4-byte register
-- Architecture : structural
-- Author: Daniel Giro, Ian Lane
--

entity 4byte_reg is
  port(

  );
end 4byte_reg;
