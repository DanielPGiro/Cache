--
-- Entity: counter_reg
-- Architecture : structural
-- Author: giropau1
-- Created On: 11/15/2014
--
library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity counter_reg is
  port (
    clk     : in  std_logic;
    rst		: in  std_logic;
    Q       : inout std_logic_vector(4 downto 0));
end counter_reg;

architecture structural of counter_reg is

component inverter
  port (
    input  : in  std_logic;
    output : out std_logic);
end component;

component dff
	port ( d   : in  std_logic;
         clk : in  std_logic;
         q   : out std_logic;
         qbar: out std_logic); 
end component;

component and2 
  port (
    input1	: in  std_logic;
	input2	: in  std_logic;
    output  : out std_logic);
end component;

component and3
  port (
    input1	: in  std_logic;
	input2	: in  std_logic;
	input3	: in  std_logic;
    output  : out std_logic);
end component;

component xor2
  port (
    input1	: in  std_logic;
	input2	: in  std_logic;
    output  : out std_logic);
end component;



for inv_0, inv_1 : inverter use entity work.inverter(structural);
for dff_0, dff_1, dff_2, dff_3, dff_4 : dff use entity work.dff(structural);
for xor2_0, xor2_1, xor2_2, xor2_3 : xor2 use entity work.xor2(structural);
for and2_0, and2_1, and2_2, and2_3, and2_4, and2_5, and2_6 : and2 use entity work.and2(structural);
for and3_0, and3_1 : and3 use entity work.and3(structural);


signal rst_bar, Q0_bar	: std_logic;
signal temp1 	: std_logic;
signal temp2	: std_logic_vector (1 downto 0);
signal temp3 	: std_logic_vector (1 downto 0);
signal temp4	: std_logic_vector (2 downto 0);
signal Q_temp, Qin	: std_logic_vector (4 downto 0);

begin

inv_0 : inverter port map (rst, rst_bar);

-- Bit 0 --
inv_1 : inverter port map (Q(0), Q0_bar);
and2_0: and2 port map (Q0_bar, rst_bar, Q_temp(0));
dff_0: dff port map (Q_temp(0), clk, Q(0));

-- Bit 1 --
xor2_0: xor2 port map (Q(0), Q(1), temp1);
and2_1: and2 port map (temp1, rst_bar, Q_temp(1));
dff_1: dff port map (Q_temp(1), clk, Q(1));

-- Bit 2 -- 
and2_2: and2 port map (Q(0), Q(1), temp2(0)); 
xor2_1: xor2 port map (Q(2), temp2(0), temp2(1));
and2_3: and2 port map (temp2(1), rst_bar, Q_temp(2));
dff_2: dff port map (Q_temp(2), clk, Q(2));

-- Bit 3 -- 
and3_0: and3 port map (Q(0), Q(1), Q(2), temp3(0));
xor2_2: xor2 port map (Q(3), temp3(0), temp3(1));
and2_4: and2 port map (temp3(1), rst_bar, Q_temp(3));
dff_3: dff port map (Q_temp(3), clk, Q(3));

-- Bit 4 --  
and3_1: and3 port map (Q(0), Q(1), Q(2), temp4(0));
and2_5: and2 port map (Q(3), temp4(0), temp4(1)); 
xor2_3: xor2 port map (Q(4), temp4(1), temp4(2));
and2_6: and2 port map (temp4(2), rst_bar, Q_temp(4));
dff_4: dff port map (Q_temp(4), clk, Q(4));

end structural;

