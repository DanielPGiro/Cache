-- Created by @(#)$CDS: vhdlin version IC23.1-64b 06/21/2023 09:20 (cpgbld16) $
-- on Mon Nov  3 12:21:32 2025


architecture structural of or7 is
begin
  output <= input1 or input2 or input3 or input4 or input5 or input6 or input7;

end structural;
