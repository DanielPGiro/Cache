--
-- Entity: negative edge triggered registers (reg)
-- Architecture : structural
-- Author: Daniel Giro, Ian Lane
--

entity reg is
  port (
    

  );
end reg;
