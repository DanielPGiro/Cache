-- Created by @(#)$CDS: vhdlin version IC23.1-64b 06/21/2023 09:20 (cpgbld16) $
-- on Mon Nov  3 12:21:32 2025


architecture structural of dff_p is

begin
  
  output: process

  begin
    wait until (clk'EVENT and clk = '1');
    q <= d;
    qbar <= not d;
  end process output;

end structural;
