--
-- Entity: negative edge triggered cache memory (cache_mem)
-- Architecture: structural
-- Author: Daniel Giro, Ian Lane

library IEEE;
library STD;
use IEEE.std_logic_1164.all;


entity current_state is
  port (
    
  );
end current_state;

architecture structural of current_state is
  component 
    port (
      
    );
  end component;

for curr_s: use entity ;

signal ;

begin


end structural;
