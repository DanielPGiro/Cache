--
-- Entity: negative edge triggered cache memory (cache_mem)
-- Architecture : structural
-- Author: Daniel Giro, Ian Lane
--

entity cache_mem is
  port (

  );
end cache_mem;

  
