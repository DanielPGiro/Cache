--
-- Entity: negative edge triggered cache memory (cache_mem)
-- Architecture: structural
-- Author: Daniel Giro, Ian Lane

library IEEE;
library STD;
use IEEE.std_logic_1164.all;


entity  is
  port (
    
  );

end cache mem;

architecture structural of current_state is
  component 
    port (
      
    );
  end component;

for cs: use entity ;

signal ;

begin


end structural;
