--
-- Entity: negative edge triggered state machine
-- Architecture : structural
-- Author: Daniel Giro, Ian Lane
--

entity state_machine is
  port( 

  );
end state_machine;
