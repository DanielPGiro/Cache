--
-- Entity: negative edge triggered ram
-- Architecture : structural
-- Author: Daniel Giro, Ian Lane
--

entity ram is
  port (
    

  );
end ram
