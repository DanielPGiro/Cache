--
-- Entity: negative edge triggered block (4-byte register)
-- Architecture : structural
-- Author: Daniel Giro, Ian Lane
-- There will be four of these in the cache, totaling 16 bytes
--

entity 4byte_reg is
  port(

  );
end 4byte_reg;
