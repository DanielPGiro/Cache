--
-- Entity: negative edge triggered hit_miss_logic
-- Architecture : structural
-- Author: Daniel Giro, Ian Lane
--

entity hit_miss_logic is
  port (

  );
end hit_miss_logic;
